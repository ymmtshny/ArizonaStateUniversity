`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:43:25 04/22/2016
// Design Name:   Project3_TestBench_byInstructor
// Module Name:   C:/Xilinx/14.7/ISE_DS/ISE/Shinya_Yamamoto/Project3_Shinya_Yamamoto/Project3_TestBench_by_Shinya_Yamamoto.v
// Project Name:  Project3_Shinya_Yamamoto
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Project3_TestBench_byInstructor
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Project3_TestBench_by_Shinya_Yamamoto;

	// Instantiate the Unit Under Test (UUT)
	Project3_TestBench_byInstructor uut (
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

