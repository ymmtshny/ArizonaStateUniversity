`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:00:34 07/05/2015
// Design Name:   Project3
// Module Name:   C:/Users/yhidalgo/Documents/ser232/Yoalli_Project3/Project3_TestBench_byInstructor.v
// Project Name:  Project3
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Project3
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Project3_TestBench_byInstructor;

	// Inputs
	reg [3:0] opCode;
	reg signed [15:0] in1;
	reg signed [15:0] in2;
	
	
	// Outputs
	wire signed [15:0] result;
	wire overflow;

	// Internal registers
	reg signed [15:0] expectedResult;
	reg expectedOverflow;
	
	// Instantiate the Unit Under Test (UUT)
	calculator uut (
		.result(result), 
		.overflow(overflow), 
		.opCode(opCode), 
		.in1(in1), 
		.in2(in2)
	);
	integer numberOfCorrectTestCases;
	integer numberOfIncorrectTestCases;
	always@(in1, in2, opCode)begin
		#25; //Allow some time to make sure result and overflow get updated in the calculator. 
		if( (result==expectedResult) & (overflow==expectedOverflow) ) begin
			numberOfCorrectTestCases = numberOfCorrectTestCases+1;
		end
		else begin 
			$display("");//The following two lines display the same, just one in binary and the other in decimal:
			$display("in1=%b in2=%b opCode=%b result= %b  expectedResult= %b     overflow=%b expectedOverflow=%b", in1, in2, opCode, result, expectedResult, overflow, expectedOverflow);
			$display("in1=%d           in2=%d           opCode=%d     result= %d            expectedResult= %d               overflow=%d  expectedOverflow=%d", in1, in2, opCode, result, expectedResult, overflow, expectedOverflow);
			numberOfIncorrectTestCases = numberOfIncorrectTestCases+1;
		end
	end
	initial begin
		// Initialize Inputs and internal registers/variables
		numberOfCorrectTestCases = 0;
		numberOfIncorrectTestCases = 0;
		opCode = 0;
		in1 = 0;
		in2 = 0;
		expectedOverflow='b0; 
		expectedResult='b0000000000000000;

		// Wait 100 ns for global reset to finish
		#100;
      $display("IMPORTANT: Make sure the Simulation lasts for at least 145000 ns, to ensure all test cases run. ");
		
		//Test opCode=0000
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0000; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000100; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011100; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001011; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110010111; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110011000; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0001100110011100; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001110; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110011000; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110011001; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001011; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100100; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100101; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100110; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110000; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110001; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100101; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100110; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100111; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110001; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b0100110011001110; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100110; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001100111; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b0110011001101000; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110010111; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110011000; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110000; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110001; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110010; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1111111111111100; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1111111111111101; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0000; expectedOverflow='b1; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110011000; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0000; expectedOverflow='b1; expectedResult='b1001100110011001; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110001; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110010; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0000; expectedOverflow='b1; expectedResult='b1011001100110011; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0000; expectedOverflow='b1; expectedResult='b1111111111111101; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0000; expectedOverflow='b1; expectedResult='b1111111111111110; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0000; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0000; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0000; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0000; expectedOverflow='b1; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0000; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0000; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0000; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0000; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0000; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0000; expectedOverflow='b1; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0000; expectedOverflow='b1; expectedResult='b0000000000000010; #100; 
		//Test opCode=0001
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100111; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001110; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001101000; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100111; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001111; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001110; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001101001; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001101000; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011010000; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001111; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b1100110011001110; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000100; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1000000000000001; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110010111; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100111; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1001100110011001; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1001100110011000; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001101000; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100111; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1001100110011100; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1001100110011010; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1001100110011001; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110000; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1011001100110001; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b1011001100110110; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1011001100110100; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1011001100110011; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0111111111111100; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b0110011001100101; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b0110011001100100; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b0100110011001011; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b0100110011001010; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1111111111111110; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1111111111111101; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0001; expectedOverflow='b0; expectedResult='b0110011001100110; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0001; expectedOverflow='b0; expectedResult='b0110011001100101; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0001; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0001; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0001; expectedOverflow='b0; expectedResult='b0100110011001011; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0001; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b1111111111111110; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0001; expectedOverflow='b1; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0001; expectedOverflow='b1; expectedResult='b0110011001100111; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0001; expectedOverflow='b1; expectedResult='b0110011001100110; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0001; expectedOverflow='b1; expectedResult='b0100110011001110; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0001; expectedOverflow='b1; expectedResult='b0100110011001101; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0001; expectedOverflow='b1; expectedResult='b0100110011001100; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0001; expectedOverflow='b1; expectedResult='b0000000000000010; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0001; expectedOverflow='b1; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0001; expectedOverflow='b1; expectedResult='b0110011001101000; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0001; expectedOverflow='b1; expectedResult='b0110011001100111; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0001; expectedOverflow='b1; expectedResult='b0100110011001111; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0001; expectedOverflow='b1; expectedResult='b0100110011001110; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0001; expectedOverflow='b1; expectedResult='b0100110011001101; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0001; expectedOverflow='b1; expectedResult='b0000000000000011; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0001; expectedOverflow='b1; expectedResult='b0000000000000010; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		//Test opCode=0010
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000000101; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0000000000001010; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0010; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000010; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111010; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1111111111111111; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b0000000000000100; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111110110; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b0111111111111011; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0010; expectedOverflow='b1; expectedResult='b1000000000000101; #100; 
		//Test opCode=0011
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0011; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000001010001111; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000010100011110; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b0000110011001100; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0011; expectedOverflow='b1; expectedResult='b1111001100110100; #100; 
		//Test opCode=0100
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010000; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010001; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010000; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010010; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010010; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010000; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010000; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010010; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110000; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010001; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010010; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110000; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010000; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001000100010000; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110000; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110000; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0100; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0100; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0100; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		//Test opCode=0101
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110000; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111100; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101011; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101010; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101101; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100111; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100110; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011000; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101000; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101001; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101110; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100100; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100101; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110000; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101011; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101000; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000110; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101010; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101001; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000111; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101101; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0010101010101110; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000110; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000111; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001010; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001011; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111100; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100111; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100100; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001010; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100110; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b0110011001100101; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001101; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001100; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b0100110011001011; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0101; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011000; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0101; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0101; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0101; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0101; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		//Test opCode=0110
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111011; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111011; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111101; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111010; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111011; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111110; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111011; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111010; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111011; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111011; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110111; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111101; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011101110111110; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110110; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110111; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011010; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110010; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110100; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000011; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011001; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0110; expectedOverflow='b0; expectedResult='b1001100110011011; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110011; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0110; expectedOverflow='b0; expectedResult='b1011001100110101; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0110; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0110; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		//Test opCode=0111
		in1='b0000000000000000; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111110; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1111111111111101; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100110; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1110011001100101; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001101; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001100; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1100110011001011; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b0111; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		//Test opCode=1000
		in1='b0000000000000000; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000010; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0000000000000011; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011010; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0001100110011011; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110100; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0011001100110101; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b0111111111111111; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b1000; expectedOverflow='b1; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000001; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b1000; expectedOverflow='b0; expectedResult='b1000000000000010; #100; 
		//Test opCode=1001
		in1='b0000000000000000; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000000; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b1111111111111111; #100; 
		in1='b0000000000000001; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000001; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000000; #100; 
		in1='b0000000000000010; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0000000000000010; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0000000000000001; #100; 
		in1='b0001100110011001; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011001; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011000; #100; 
		in1='b0001100110011010; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0001100110011010; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0001100110011001; #100; 
		in1='b0011001100110010; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110010; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110001; #100; 
		in1='b0011001100110011; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110011; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110010; #100; 
		in1='b0011001100110100; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0011001100110100; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0011001100110011; #100; 
		in1='b0111111111111110; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111110; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111101; #100; 
		in1='b0111111111111111; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b0111111111111111; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b0111111111111110; #100; 
		in1='b1000000000000000; in2='b0000000000000000; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0000000000000001; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0000000000000010; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0001100110011001; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0001100110011010; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0011001100110010; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0011001100110011; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0011001100110100; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0111111111111110; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b0111111111111111; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b1000000000000000; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000000; in2='b1000000000000001; opCode='b1001; expectedOverflow='b1; expectedResult='b0111111111111111; #100; 
		in1='b1000000000000001; in2='b0000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0000000000000010; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0001100110011001; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0001100110011010; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0011001100110010; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0011001100110011; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0011001100110100; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0111111111111110; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b0111111111111111; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b1000000000000000; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		in1='b1000000000000001; in2='b1000000000000001; opCode='b1001; expectedOverflow='b0; expectedResult='b1000000000000000; #100; 
		
		
		#100;		
		$display("Number of correct test cases: %d",numberOfCorrectTestCases);
		$display("Number of incorrect test cases: %d  <- Make sure this number is zero",numberOfIncorrectTestCases);
		#100;
		
	end 
endmodule